module top(
    input a,
    input b,
    output f
);

    wire aa;
    assign aa = ~aa;
endmodule
